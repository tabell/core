`timescale 1ns/ps

module core(
	input clk;

)
subcomponent alu1 (

	)
endmodule;