`timescale 1ns / 1ps

module core(
	input clk,
	input rst,
	input clk_en
);

wire [31:0] icache_read_data;
reg [5:0] icache_read_addr;
wire icache_data_ready;
reg icache_clk_en;

l1_cache icache(
	.read_data(icache_read_data),
	.read_addr(pc[5:0]),
	.data_ready(icache_data_ready),
	.clk(clk),
	.clk_en(icache_clk_en),
	.rst(rst)
	);

wire [31:0] alu_operand_a;
reg [31:0] alu_operand_b_mux;
reg [5:0] alu_func_mux;
wire [31:0] alu_result;
reg alu_clk_en;

alu alu1(
	.operand_a(alu_operand_a),
	.operand_b(alu_operand_b_mux),
	.result(alu_result),
	.func(alu_func_mux),
	.clk(clk),
	.clk_en(alu_clk_en)
	);

wire [31:0] regfile_read_data_a;
wire [31:0] regfile_read_data_b;
reg [31:0] regfile_write_data;
reg [4:0] regfile_write_addr;
reg regfile_write_enable;

regfile regfile(
    .read_data_a(alu_operand_a),
    .read_data_b(regfile_read_data_b),
    .write_data(regfile_write_data),
    .read_addr_a(icache_read_data[25:21]),
    .read_addr_b(icache_read_data[20:16]),
    .write_addr(regfile_write_addr),
    .write_enable(regfile_write_enable),
    .clk(clk),
    .rst(rst)
    );

	wire clk;
	reg tmp=0;

	reg [15:0] pc; // program counter
	reg [15:0] n_pc; // next program counter


	reg [5:0]  exec_opcode;
	reg [15:0] exec_imm;
	reg [4:0]  exec_reg_t;
	reg [4:0]  exec_reg_d;
	reg [5:0]  exec_func;

	reg [5:0]  wb_opcode;
	reg [15:0] wb_imm;
	reg [4:0]  wb_reg_t;


	reg alu_operand_b_mux_sel;
	reg alu_func_mux_sel;


always @(posedge clk or posedge rst) begin
	if(rst) begin
		// reset PC
		pc <= 0; // start address 10 so maybe interrupts later?
		n_pc <= 10;

		// clock enables
		icache_clk_en <= 0;
		alu_clk_en <= 0;

	end else if(clk_en) begin
		// on every cycle
		// set new PC
		if (decode_opcode == 2)
			n_pc <= n_pc + decode_sign_imm[15:0];
		else
			n_pc <= n_pc + 1;
		pc <= n_pc;

		// clock enables
		icache_clk_en <= 1;
		alu_clk_en <= 1;

		// fetch stage
		// icache_read_addr <= n_pc[5:0];

		// decode

		// execute
		regfile_write_enable <= 0;
		regfile_write_addr <= 5'hZ;

		exec_opcode <= decode_opcode;
		exec_reg_t <= decode_reg_t;
		exec_reg_d <= decode_reg_d;
		exec_imm <= decode_imm;
		exec_func <= decode_func;

		// writeback
		wb_imm <= exec_imm;
		wb_opcode <= exec_opcode;
		wb_reg_t <= exec_reg_t;
		
		if (exec_opcode == 15) begin // load immediate hi
			regfile_write_addr <= exec_reg_t;
			regfile_write_enable <= 1;
			regfile_write_data <= exec_imm;
			// assign regfile_write_data = {wb_imm,{16{1'b0}}};
		end else if (exec_opcode == 0) begin
			if (exec_reg_d == 0)
				regfile_write_enable <= 0;
			else begin
				regfile_write_enable <= 1;
				regfile_write_addr <= exec_reg_d;
				regfile_write_data <= alu_result;
			end
		end else if (exec_opcode == 8) begin // add immediate
			regfile_write_enable <= 1;
			regfile_write_addr <= exec_reg_t;
			regfile_write_data <= alu_result;
		end

		// switches ALU input b betwen regfile output and
		// decoded immediate value
		if (decode_opcode == 8)
			alu_operand_b_mux_sel <= 0;
		else
			alu_operand_b_mux_sel <= 1;
		// switches alu func input between decoded
		// func and decoded opcode

	end
end

wire [25:0] decode_full_imm = icache_read_data[25:0];
wire [5:0] decode_opcode = icache_read_data[31:26];
wire [4:0] decode_reg_s = icache_read_data[25:21]; // source a
wire [4:0] decode_reg_t = icache_read_data[20:16]; // source b
wire [4:0] decode_reg_d = icache_read_data[15:11]; // dest
wire [4:0] decode_shamt = icache_read_data[10:6]; // shift amount
wire [5:0] decode_func = icache_read_data[5:0]; // alu function
wire [15:0] decode_imm = icache_read_data[15:0];
wire [31:0] decode_sign_imm = {{6{icache_read_data[25]}},icache_read_data[25:0]};

// alu_operand_b = alu_operand_b_mux_sel ? read_data_b : decode_imm;
always @(*) begin
	case (decode_opcode)
		8 : alu_operand_b_mux <= decode_imm;
		default : alu_operand_b_mux <= regfile_read_data_b;
	endcase




	case (decode_opcode)
		0 :	alu_func_mux <= decode_func;
		default : alu_func_mux <= decode_opcode;
	endcase




end
    
endmodule