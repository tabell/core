`define func_add 0'b100000
`define func_addu 0'b100001
`define func_addi 0'b001000
`define func_addiu 0'b001001
`define func_and 0'b100100
`define func_andi 0'b001100
`define func_div 0'b011010
`define func_divu 0'b011011
`define func_mult 0'b011000
`define func_multu 0'b011001
`define func_nor 0'b100111
`define func_or 0'b100101
`define func_ori 0'b001101
`define func_sll 0'b000000
`define func_sllv 0'b000100
`define func_sra 0'b000011
`define func_srav 0'b000111
`define func_srl 0'b000010
`define func_srlv 0'b000110
`define func_sub 0'b100010
`define func_subu 0'b100011
`define func_xor 0'b100110
`define func_xori 0'b001110